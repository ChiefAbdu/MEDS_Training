// new logic
